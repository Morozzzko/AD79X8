module TestBench();
endmodule
