module ADC(in, out, sclk, reset);
endmodule
